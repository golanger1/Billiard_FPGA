// (c) Technion IIT, Department of Electrical Engineering 2020 

// Implements a slow clock as an one-second counter
// Turbo input sets output 10 times faster
// Updated by Mor Dahan - January 2022

 
 module one_sec_counter      	
	(
   // Input, Output Ports
	input  logic clk, 
	input  logic resetN, 
	input  logic turbo,
	output logic one_sec
   );
	
	int oneSecCount ;
	int sec ;		 // gets either one seccond or Turbo top value

// counter limit setting 
	
//       ----------------------------------------------	
	localparam oneSecVal = 26'd25_000_000; // for DE10 board un-comment this line 
//	localparam oneSecVal = 26'd50_000_000; // for DE10 board un-comment this line 
//	localparam oneSecVal = 26'd20; // for quartus simulation un-comment this line 
//       ----------------------------------------------	
	
	assign  sec = turbo ? oneSecVal/10 : oneSecVal;  // it is legal to devide by 10, as it is done by the complier not by logic (actual transistors) 


	
   always_ff @( posedge clk or negedge resetN )
   begin
	
		// asynchronous reset
		if ( !resetN ) 
			begin
				one_sec <= 1'b0;
				oneSecCount <= 0;
			end // if reset
		
		// executed once every clock 	
		else 
			begin
				if (oneSecCount >= sec) 
					begin
						oneSecCount <= 0;
						one_sec		<= 1'b1;
					end
				else 
					begin
						oneSecCount <= oneSecCount + 1;
						one_sec		<= 1'b0;
					end
			end // else clk
		
	end // always
endmodule